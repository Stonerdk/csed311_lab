module sign_extender(in, out);
input reg[7:0] in;
output reg[15:0] out;
begin
    // TODO
end